# asynchronous-fifo
<br>
AUthor Mihir Kalaariya (changed)
AUthor Mihir Kalaariya (changed)
AUthor Mihir Kalaariya (changed)
AUthor Mihir Kalaariya (changed)
AUthor Mihir Kalaariya (changed)
